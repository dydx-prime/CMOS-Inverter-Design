magic
tech sky130A
timestamp 1752193593
<< nwell >>
rect -110 30 185 320
<< nmos >>
rect 35 -145 50 -45
<< pmos >>
rect 35 60 50 260
<< ndiff >>
rect -15 -65 35 -45
rect -15 -120 -5 -65
rect 15 -120 35 -65
rect -15 -145 35 -120
rect 50 -65 100 -45
rect 50 -120 70 -65
rect 90 -120 100 -65
rect 50 -145 100 -120
<< pdiff >>
rect -15 205 35 260
rect -15 150 -5 205
rect 15 150 35 205
rect -15 60 35 150
rect 50 205 100 260
rect 50 150 70 205
rect 90 150 100 205
rect 50 60 100 150
<< ndiffc >>
rect -5 -120 15 -65
rect 70 -120 90 -65
<< pdiffc >>
rect -5 150 15 205
rect 70 150 90 205
<< poly >>
rect 35 260 50 280
rect 35 35 50 60
rect -10 25 50 35
rect -10 5 0 25
rect 20 5 50 25
rect -10 -5 50 5
rect 35 -45 50 -5
rect 35 -160 50 -145
<< polycont >>
rect 0 5 20 25
<< locali >>
rect -40 285 30 305
rect 55 285 120 305
rect -15 205 20 285
rect -15 150 -5 205
rect 15 150 20 205
rect -15 60 20 150
rect 65 205 100 260
rect 65 150 70 205
rect 90 150 100 205
rect -10 25 30 35
rect -10 5 0 25
rect 20 5 30 25
rect -10 -5 30 5
rect -15 -65 20 -45
rect -15 -120 -5 -65
rect 15 -120 20 -65
rect -15 -180 20 -120
rect 65 -65 100 150
rect 65 -120 70 -65
rect 90 -120 100 -65
rect 65 -145 100 -120
rect -40 -200 30 -180
rect 55 -200 120 -180
<< viali >>
rect -65 285 -40 305
rect 30 285 55 305
rect 120 285 145 305
rect -65 -200 -40 -180
rect 30 -200 55 -180
rect 120 -200 145 -180
<< metal1 >>
rect -80 305 155 310
rect -80 285 -65 305
rect -40 285 30 305
rect 55 285 120 305
rect 145 285 155 305
rect -80 280 155 285
rect -75 -180 160 -175
rect -75 -200 -65 -180
rect -40 -200 30 -180
rect 55 -200 120 -180
rect 145 -200 160 -180
rect -75 -205 160 -200
<< labels >>
rlabel viali 30 285 55 305 1 Vdd
rlabel polycont 0 5 20 25 1 Vin
rlabel locali 65 0 100 30 1 Vout
rlabel viali 30 -200 55 -180 1 gnd
rlabel nwell -110 30 185 320 1 Vdd
<< end >>
