magic
tech sky130A
timestamp 1751245013
<< nwell >>
rect -50 -50 250 355
<< nmos >>
rect 90 -200 105 -100
<< pmos >>
rect 90 0 105 200
<< ndiff >>
rect 45 -110 90 -100
rect 45 -190 55 -110
rect 75 -190 90 -110
rect 45 -200 90 -190
rect 105 -110 150 -100
rect 105 -190 120 -110
rect 140 -190 150 -110
rect 105 -200 150 -190
<< pdiff >>
rect 40 190 90 200
rect 40 10 50 190
rect 75 10 90 190
rect 40 0 90 10
rect 105 190 155 200
rect 105 10 120 190
rect 145 10 155 190
rect 105 0 155 10
<< ndiffc >>
rect 55 -190 75 -110
rect 120 -190 140 -110
<< pdiffc >>
rect 50 10 75 190
rect 120 10 145 190
<< psubdiff >>
rect 45 -245 150 -230
rect 45 -265 60 -245
rect 135 -265 150 -245
rect 45 -280 150 -265
<< nsubdiff >>
rect 25 305 175 320
rect 25 275 40 305
rect 160 275 175 305
rect 25 260 175 275
<< psubdiffcont >>
rect 60 -265 135 -245
<< nsubdiffcont >>
rect 40 275 160 305
<< poly >>
rect 90 200 105 250
rect 90 -100 105 0
rect 90 -215 105 -200
<< locali >>
rect 25 305 175 320
rect 25 275 40 305
rect 160 275 175 305
rect 25 260 175 275
rect 40 190 85 200
rect 40 10 50 190
rect 75 10 85 190
rect 40 0 85 10
rect 110 190 155 200
rect 110 10 120 190
rect 145 10 155 190
rect 110 0 155 10
rect 45 -110 85 -100
rect 45 -190 55 -110
rect 75 -190 85 -110
rect 45 -200 85 -190
rect 110 -110 150 -100
rect 110 -190 120 -110
rect 140 -190 150 -110
rect 110 -200 150 -190
rect 45 -245 150 -230
rect 45 -265 60 -245
rect 135 -265 150 -245
rect 45 -280 150 -265
<< end >>
