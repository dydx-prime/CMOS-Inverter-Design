** sch_path: /home/prime/CMOS-Inverter-Design/schematics/inv.sch
**.subckt inv
Vdd Vdd gnd 1.8
Vin Vin gnd PULSE(0 1.8 0 .3n .3n 3n 6.6n 5)
C1 Vout net1 0p m=1
X0 Vout Vin gnd gnd sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
**** begin user architecture code

.lib /home/prime/vlsi_/open_pdks/sources/sky130_fd_pr/models/sky130.lib.spice tt
.dc Vin 0 2 1m
.tran .02n 10n
.save all
.end

**** end user architecture code
**.ends
.GLOBAL gnd
.end

